module runtime

import types